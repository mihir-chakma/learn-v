module main

fn main() {
	println('Hello World!')
}

// this is a single comment 
/*
   Multiline comment
*/
